`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:29:59 04/20/2019 
// Design Name: 
// Module Name:    trab1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module trab1(
    input count,
    input up_down,
    input load,
    input [3:0] load_input,
    input reset,
    input clk
    );


endmodule
